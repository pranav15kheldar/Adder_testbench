interface inf_adder();
    logic clk;
    logic a;
    logic b;
    logic c;
    logic sum;
    logic carry;
endinterface