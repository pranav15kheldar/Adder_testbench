class transaction;
    rand logic a;
    rand logic b;
    rand logic c;
    logic sum;
    logic carry;
endclass