package adder;
    `include "transaction.sv"
    `include "generator.sv"
    `include "driver.sv"
    `include "enviroment.sv"
    `include "test.sv"
endpackage